// ===============================================================
// vu_meter_6led.sv
// 6-LED VU-meter for 24-bit PCM audio samples
// Consumes samples from ram_logic via ready/valid handshake
// ===============================================================
module vu_meter_6led #(
  // Leaky integrator parameters
  parameter int DECAY_SHIFT    = 14,        // Decay rate: higher = slower decay (12-16 recommended)
  parameter int SCALE_SHIFT    = 2,         // Sensitivity: higher = less sensitive (0-4 recommended)

  // LED threshold levels (32-bit to match level_q width)
  parameter int unsigned TH1   = 32'd500,   // LED 1 threshold
  parameter int unsigned TH2   = 32'd2000,  // LED 2 threshold
  parameter int unsigned TH3   = 32'd6000,  // LED 3 threshold
  parameter int unsigned TH4   = 32'd15000, // LED 4 threshold
  parameter int unsigned TH5   = 32'd35000, // LED 5 threshold
  parameter int unsigned TH6   = 32'd70000, // LED 6 threshold

  // LED refresh rate: ~50 Hz at 27 MHz clock
  parameter int LED_DIV        = 540000     // 27e6 / 540000 = 50 Hz
)(
  input  logic               clk_i,             // System clock (27 MHz)
  input  logic               rst_ni,            // Active-low reset

  // RAM consumer interface (ready/valid handshake)
  input  logic signed [23:0] ram_read_data_i,   // Sample data from RAM
  input  logic               ram_read_valid_i,  // Valid signal from RAM
  output logic               ram_read_ready_o,  // Ready signal to RAM

  input  logic               ram_buffer_ready_i, // Buffer ready indicator (optional monitoring)

  // LED outputs
  output logic [5:0]         leds_o             // LED control signals
);

  //==========================================================================
  // Internal signals
  //==========================================================================

  // Processing state machine
  typedef enum logic [1:0] {
    IDLE,       // Ready to accept new sample
    COMPUTE,    // Computing magnitude and updating level
    SETTLE      // Allowing computation to settle
  } state_t;

  state_t state_q, state_d;

  // Sample processing
  logic signed [23:0] sample_q;          // Registered input sample
  logic        [23:0] magnitude;         // Absolute value of sample
  logic               sample_accepted;   // Handshake occurred

  // Level tracking
  logic        [31:0] level_q, level_d;  // Leaky integrator output

  // LED update control
  logic [$clog2(LED_DIV)-1:0] refresh_counter_q;
  logic                        led_update_tick;

  //==========================================================================
  // Ready/valid handshake
  //==========================================================================
  assign sample_accepted = ram_read_valid_i && ram_read_ready_o;
  assign ram_read_ready_o = (state_q == IDLE);

  //==========================================================================
  // Magnitude calculation (absolute value)
  //==========================================================================
  always_comb begin
    magnitude = sample_q[23] ? (~sample_q + 24'b1) : sample_q;
  end

  //==========================================================================
  // State machine for sample processing
  //==========================================================================
  always_comb begin
    // Default: maintain state
    state_d = state_q;
    level_d = level_q;

    case (state_q)
      IDLE: begin
        if (sample_accepted) begin
          // Sample handshake occurred, start processing
          state_d = COMPUTE;
        end
      end

      COMPUTE: begin
        // Update leaky integrator: decay old level, add new scaled magnitude
        level_d = level_q - (level_q >> DECAY_SHIFT) + (magnitude >> SCALE_SHIFT);
        state_d = SETTLE;
      end

      SETTLE: begin
        // Allow computation to settle, then return to idle
        state_d = IDLE;
      end

      default: state_d = IDLE;
    endcase
  end

  // State and level register
  always_ff @(posedge clk_i) begin
    if (!rst_ni) begin
      state_q  <= IDLE;
      level_q  <= 32'd0;
      sample_q <= 24'd0;
    end else begin
      state_q <= state_d;
      level_q <= level_d;
      if (sample_accepted) begin
        sample_q <= ram_read_data_i;
      end
    end
  end

  //==========================================================================
  // LED refresh rate divider (~50 Hz to prevent flicker)
  //==========================================================================
  always_ff @(posedge clk_i) begin
    if (!rst_ni) begin
      refresh_counter_q <= '0;
      led_update_tick   <= 1'b0;
    end else begin
      if (refresh_counter_q == LED_DIV - 1) begin
        refresh_counter_q <= '0;
        led_update_tick   <= 1'b1;
      end else begin
        refresh_counter_q <= refresh_counter_q + 1'b1;
        led_update_tick   <= 1'b0;
      end
    end
  end

  //==========================================================================
  // LED threshold comparison and output
  //==========================================================================
  logic [5:0] leds_d;

  always_comb begin
    leds_d[0] = (level_q >= TH1);
    leds_d[1] = (level_q >= TH2);
    leds_d[2] = (level_q >= TH3);
    leds_d[3] = (level_q >= TH4);
    leds_d[4] = (level_q >= TH5);
    leds_d[5] = (level_q >= TH6);
  end

  // Update LED outputs only on refresh tick to reduce flicker
  always_ff @(posedge clk_i) begin
    if (!rst_ni) begin
      leds_o <= 6'b0;
    end else if (led_update_tick) begin
      leds_o <= leds_d;
    end
  end

endmodule
