// ============================================================================
// fpga_template_pkg.sv
// Package for FPGA template project - type definitions and constants
// ============================================================================

package fpga_template_pkg;

  // Add type definitions and constants here as needed
  // Currently empty - reserved for future use

endpackage : fpga_template_pkg
