// ============================================================================
// fft_twiddle_256 - Twiddle Factor ROM for 256-Point FFT
// ============================================================================
// Precomputed twiddle factors (complex exponentials) for FFT
//
// Twiddle factors: W_N^k = e^(-j*2*pi*k/N) = cos(2πk/N) - j*sin(2πk/N)
// Format: Q1.17 (18-bit signed fixed-point, 17 fractional bits)
// Range: -1.0 to +0.999992370 represented as -131072 to +131071
// ============================================================================

module fft_twiddle_256 #(
    parameter int DATA_WIDTH = 18
) (
    input  logic                    clk_i,
    input  logic [7:0]              addr_i,     // Twiddle factor index (0-255)
    output logic signed [DATA_WIDTH-1:0] cos_o, // Real part (cosine)
    output logic signed [DATA_WIDTH-1:0] sin_o  // Imaginary part (-sine for FFT)
);

    // Synchronous ROM
    always_ff @(posedge clk_i) begin
        case (addr_i)
            8'd0:   begin cos_o = 18'sd131071;  sin_o = 18'sd0; end
            8'd1:   begin cos_o = 18'sd131032;  sin_o = -18'sd3216; end
            8'd2:   begin cos_o = 18'sd130914;  sin_o = -18'sd6431; end
            8'd3:   begin cos_o = 18'sd130716;  sin_o = -18'sd9642; end
            8'd4:   begin cos_o = 18'sd130440;  sin_o = -18'sd12847; end
            8'd5:   begin cos_o = 18'sd130086;  sin_o = -18'sd16044; end
            8'd6:   begin cos_o = 18'sd129653;  sin_o = -18'sd19232; end
            8'd7:   begin cos_o = 18'sd129142;  sin_o = -18'sd22408; end
            8'd8:   begin cos_o = 18'sd128553;  sin_o = -18'sd25570; end
            8'd9:   begin cos_o = 18'sd127887;  sin_o = -18'sd28718; end
            8'd10:   begin cos_o = 18'sd127143;  sin_o = -18'sd31847; end
            8'd11:   begin cos_o = 18'sd126324;  sin_o = -18'sd34958; end
            8'd12:   begin cos_o = 18'sd125428;  sin_o = -18'sd38048; end
            8'd13:   begin cos_o = 18'sd124456;  sin_o = -18'sd41114; end
            8'd14:   begin cos_o = 18'sd123410;  sin_o = -18'sd44156; end
            8'd15:   begin cos_o = 18'sd122289;  sin_o = -18'sd47172; end
            8'd16:   begin cos_o = 18'sd121094;  sin_o = -18'sd50159; end
            8'd17:   begin cos_o = 18'sd119827;  sin_o = -18'sd53115; end
            8'd18:   begin cos_o = 18'sd118487;  sin_o = -18'sd56040; end
            8'd19:   begin cos_o = 18'sd117076;  sin_o = -18'sd58931; end
            8'd20:   begin cos_o = 18'sd115595;  sin_o = -18'sd61786; end
            8'd21:   begin cos_o = 18'sd114044;  sin_o = -18'sd64605; end
            8'd22:   begin cos_o = 18'sd112424;  sin_o = -18'sd67384; end
            8'd23:   begin cos_o = 18'sd110736;  sin_o = -18'sd70123; end
            8'd24:   begin cos_o = 18'sd108982;  sin_o = -18'sd72819; end
            8'd25:   begin cos_o = 18'sd107162;  sin_o = -18'sd75472; end
            8'd26:   begin cos_o = 18'sd105278;  sin_o = -18'sd78079; end
            8'd27:   begin cos_o = 18'sd103330;  sin_o = -18'sd80639; end
            8'd28:   begin cos_o = 18'sd101320;  sin_o = -18'sd83151; end
            8'd29:   begin cos_o = 18'sd99248;  sin_o = -18'sd85612; end
            8'd30:   begin cos_o = 18'sd97117;  sin_o = -18'sd88022; end
            8'd31:   begin cos_o = 18'sd94928;  sin_o = -18'sd90379; end
            8'd32:   begin cos_o = 18'sd92681;  sin_o = -18'sd92681; end
            8'd33:   begin cos_o = 18'sd90379;  sin_o = -18'sd94928; end
            8'd34:   begin cos_o = 18'sd88022;  sin_o = -18'sd97117; end
            8'd35:   begin cos_o = 18'sd85612;  sin_o = -18'sd99248; end
            8'd36:   begin cos_o = 18'sd83151;  sin_o = -18'sd101320; end
            8'd37:   begin cos_o = 18'sd80639;  sin_o = -18'sd103330; end
            8'd38:   begin cos_o = 18'sd78079;  sin_o = -18'sd105278; end
            8'd39:   begin cos_o = 18'sd75472;  sin_o = -18'sd107162; end
            8'd40:   begin cos_o = 18'sd72819;  sin_o = -18'sd108982; end
            8'd41:   begin cos_o = 18'sd70123;  sin_o = -18'sd110736; end
            8'd42:   begin cos_o = 18'sd67384;  sin_o = -18'sd112424; end
            8'd43:   begin cos_o = 18'sd64605;  sin_o = -18'sd114044; end
            8'd44:   begin cos_o = 18'sd61786;  sin_o = -18'sd115595; end
            8'd45:   begin cos_o = 18'sd58931;  sin_o = -18'sd117076; end
            8'd46:   begin cos_o = 18'sd56040;  sin_o = -18'sd118487; end
            8'd47:   begin cos_o = 18'sd53115;  sin_o = -18'sd119827; end
            8'd48:   begin cos_o = 18'sd50159;  sin_o = -18'sd121094; end
            8'd49:   begin cos_o = 18'sd47172;  sin_o = -18'sd122289; end
            8'd50:   begin cos_o = 18'sd44156;  sin_o = -18'sd123410; end
            8'd51:   begin cos_o = 18'sd41114;  sin_o = -18'sd124456; end
            8'd52:   begin cos_o = 18'sd38048;  sin_o = -18'sd125428; end
            8'd53:   begin cos_o = 18'sd34958;  sin_o = -18'sd126324; end
            8'd54:   begin cos_o = 18'sd31847;  sin_o = -18'sd127143; end
            8'd55:   begin cos_o = 18'sd28718;  sin_o = -18'sd127887; end
            8'd56:   begin cos_o = 18'sd25570;  sin_o = -18'sd128553; end
            8'd57:   begin cos_o = 18'sd22408;  sin_o = -18'sd129142; end
            8'd58:   begin cos_o = 18'sd19232;  sin_o = -18'sd129653; end
            8'd59:   begin cos_o = 18'sd16044;  sin_o = -18'sd130086; end
            8'd60:   begin cos_o = 18'sd12847;  sin_o = -18'sd130440; end
            8'd61:   begin cos_o = 18'sd9642;  sin_o = -18'sd130716; end
            8'd62:   begin cos_o = 18'sd6431;  sin_o = -18'sd130914; end
            8'd63:   begin cos_o = 18'sd3216;  sin_o = -18'sd131032; end
            8'd64:   begin cos_o = 18'sd0;  sin_o = -18'sd131072; end
            8'd65:   begin cos_o = -18'sd3216;  sin_o = -18'sd131032; end
            8'd66:   begin cos_o = -18'sd6431;  sin_o = -18'sd130914; end
            8'd67:   begin cos_o = -18'sd9642;  sin_o = -18'sd130716; end
            8'd68:   begin cos_o = -18'sd12847;  sin_o = -18'sd130440; end
            8'd69:   begin cos_o = -18'sd16044;  sin_o = -18'sd130086; end
            8'd70:   begin cos_o = -18'sd19232;  sin_o = -18'sd129653; end
            8'd71:   begin cos_o = -18'sd22408;  sin_o = -18'sd129142; end
            8'd72:   begin cos_o = -18'sd25570;  sin_o = -18'sd128553; end
            8'd73:   begin cos_o = -18'sd28718;  sin_o = -18'sd127887; end
            8'd74:   begin cos_o = -18'sd31847;  sin_o = -18'sd127143; end
            8'd75:   begin cos_o = -18'sd34958;  sin_o = -18'sd126324; end
            8'd76:   begin cos_o = -18'sd38048;  sin_o = -18'sd125428; end
            8'd77:   begin cos_o = -18'sd41114;  sin_o = -18'sd124456; end
            8'd78:   begin cos_o = -18'sd44156;  sin_o = -18'sd123410; end
            8'd79:   begin cos_o = -18'sd47172;  sin_o = -18'sd122289; end
            8'd80:   begin cos_o = -18'sd50159;  sin_o = -18'sd121094; end
            8'd81:   begin cos_o = -18'sd53115;  sin_o = -18'sd119827; end
            8'd82:   begin cos_o = -18'sd56040;  sin_o = -18'sd118487; end
            8'd83:   begin cos_o = -18'sd58931;  sin_o = -18'sd117076; end
            8'd84:   begin cos_o = -18'sd61786;  sin_o = -18'sd115595; end
            8'd85:   begin cos_o = -18'sd64605;  sin_o = -18'sd114044; end
            8'd86:   begin cos_o = -18'sd67384;  sin_o = -18'sd112424; end
            8'd87:   begin cos_o = -18'sd70123;  sin_o = -18'sd110736; end
            8'd88:   begin cos_o = -18'sd72819;  sin_o = -18'sd108982; end
            8'd89:   begin cos_o = -18'sd75472;  sin_o = -18'sd107162; end
            8'd90:   begin cos_o = -18'sd78079;  sin_o = -18'sd105278; end
            8'd91:   begin cos_o = -18'sd80639;  sin_o = -18'sd103330; end
            8'd92:   begin cos_o = -18'sd83151;  sin_o = -18'sd101320; end
            8'd93:   begin cos_o = -18'sd85612;  sin_o = -18'sd99248; end
            8'd94:   begin cos_o = -18'sd88022;  sin_o = -18'sd97117; end
            8'd95:   begin cos_o = -18'sd90379;  sin_o = -18'sd94928; end
            8'd96:   begin cos_o = -18'sd92681;  sin_o = -18'sd92681; end
            8'd97:   begin cos_o = -18'sd94928;  sin_o = -18'sd90379; end
            8'd98:   begin cos_o = -18'sd97117;  sin_o = -18'sd88022; end
            8'd99:   begin cos_o = -18'sd99248;  sin_o = -18'sd85612; end
            8'd100:   begin cos_o = -18'sd101320;  sin_o = -18'sd83151; end
            8'd101:   begin cos_o = -18'sd103330;  sin_o = -18'sd80639; end
            8'd102:   begin cos_o = -18'sd105278;  sin_o = -18'sd78079; end
            8'd103:   begin cos_o = -18'sd107162;  sin_o = -18'sd75472; end
            8'd104:   begin cos_o = -18'sd108982;  sin_o = -18'sd72819; end
            8'd105:   begin cos_o = -18'sd110736;  sin_o = -18'sd70123; end
            8'd106:   begin cos_o = -18'sd112424;  sin_o = -18'sd67384; end
            8'd107:   begin cos_o = -18'sd114044;  sin_o = -18'sd64605; end
            8'd108:   begin cos_o = -18'sd115595;  sin_o = -18'sd61786; end
            8'd109:   begin cos_o = -18'sd117076;  sin_o = -18'sd58931; end
            8'd110:   begin cos_o = -18'sd118487;  sin_o = -18'sd56040; end
            8'd111:   begin cos_o = -18'sd119827;  sin_o = -18'sd53115; end
            8'd112:   begin cos_o = -18'sd121094;  sin_o = -18'sd50159; end
            8'd113:   begin cos_o = -18'sd122289;  sin_o = -18'sd47172; end
            8'd114:   begin cos_o = -18'sd123410;  sin_o = -18'sd44156; end
            8'd115:   begin cos_o = -18'sd124456;  sin_o = -18'sd41114; end
            8'd116:   begin cos_o = -18'sd125428;  sin_o = -18'sd38048; end
            8'd117:   begin cos_o = -18'sd126324;  sin_o = -18'sd34958; end
            8'd118:   begin cos_o = -18'sd127143;  sin_o = -18'sd31847; end
            8'd119:   begin cos_o = -18'sd127887;  sin_o = -18'sd28718; end
            8'd120:   begin cos_o = -18'sd128553;  sin_o = -18'sd25570; end
            8'd121:   begin cos_o = -18'sd129142;  sin_o = -18'sd22408; end
            8'd122:   begin cos_o = -18'sd129653;  sin_o = -18'sd19232; end
            8'd123:   begin cos_o = -18'sd130086;  sin_o = -18'sd16044; end
            8'd124:   begin cos_o = -18'sd130440;  sin_o = -18'sd12847; end
            8'd125:   begin cos_o = -18'sd130716;  sin_o = -18'sd9642; end
            8'd126:   begin cos_o = -18'sd130914;  sin_o = -18'sd6431; end
            8'd127:   begin cos_o = -18'sd131032;  sin_o = -18'sd3216; end
            8'd128:   begin cos_o = -18'sd131072;  sin_o = 18'sd0; end
            8'd129:   begin cos_o = -18'sd131032;  sin_o = 18'sd3216; end
            8'd130:   begin cos_o = -18'sd130914;  sin_o = 18'sd6431; end
            8'd131:   begin cos_o = -18'sd130716;  sin_o = 18'sd9642; end
            8'd132:   begin cos_o = -18'sd130440;  sin_o = 18'sd12847; end
            8'd133:   begin cos_o = -18'sd130086;  sin_o = 18'sd16044; end
            8'd134:   begin cos_o = -18'sd129653;  sin_o = 18'sd19232; end
            8'd135:   begin cos_o = -18'sd129142;  sin_o = 18'sd22408; end
            8'd136:   begin cos_o = -18'sd128553;  sin_o = 18'sd25570; end
            8'd137:   begin cos_o = -18'sd127887;  sin_o = 18'sd28718; end
            8'd138:   begin cos_o = -18'sd127143;  sin_o = 18'sd31847; end
            8'd139:   begin cos_o = -18'sd126324;  sin_o = 18'sd34958; end
            8'd140:   begin cos_o = -18'sd125428;  sin_o = 18'sd38048; end
            8'd141:   begin cos_o = -18'sd124456;  sin_o = 18'sd41114; end
            8'd142:   begin cos_o = -18'sd123410;  sin_o = 18'sd44156; end
            8'd143:   begin cos_o = -18'sd122289;  sin_o = 18'sd47172; end
            8'd144:   begin cos_o = -18'sd121094;  sin_o = 18'sd50159; end
            8'd145:   begin cos_o = -18'sd119827;  sin_o = 18'sd53115; end
            8'd146:   begin cos_o = -18'sd118487;  sin_o = 18'sd56040; end
            8'd147:   begin cos_o = -18'sd117076;  sin_o = 18'sd58931; end
            8'd148:   begin cos_o = -18'sd115595;  sin_o = 18'sd61786; end
            8'd149:   begin cos_o = -18'sd114044;  sin_o = 18'sd64605; end
            8'd150:   begin cos_o = -18'sd112424;  sin_o = 18'sd67384; end
            8'd151:   begin cos_o = -18'sd110736;  sin_o = 18'sd70123; end
            8'd152:   begin cos_o = -18'sd108982;  sin_o = 18'sd72819; end
            8'd153:   begin cos_o = -18'sd107162;  sin_o = 18'sd75472; end
            8'd154:   begin cos_o = -18'sd105278;  sin_o = 18'sd78079; end
            8'd155:   begin cos_o = -18'sd103330;  sin_o = 18'sd80639; end
            8'd156:   begin cos_o = -18'sd101320;  sin_o = 18'sd83151; end
            8'd157:   begin cos_o = -18'sd99248;  sin_o = 18'sd85612; end
            8'd158:   begin cos_o = -18'sd97117;  sin_o = 18'sd88022; end
            8'd159:   begin cos_o = -18'sd94928;  sin_o = 18'sd90379; end
            8'd160:   begin cos_o = -18'sd92681;  sin_o = 18'sd92681; end
            8'd161:   begin cos_o = -18'sd90379;  sin_o = 18'sd94928; end
            8'd162:   begin cos_o = -18'sd88022;  sin_o = 18'sd97117; end
            8'd163:   begin cos_o = -18'sd85612;  sin_o = 18'sd99248; end
            8'd164:   begin cos_o = -18'sd83151;  sin_o = 18'sd101320; end
            8'd165:   begin cos_o = -18'sd80639;  sin_o = 18'sd103330; end
            8'd166:   begin cos_o = -18'sd78079;  sin_o = 18'sd105278; end
            8'd167:   begin cos_o = -18'sd75472;  sin_o = 18'sd107162; end
            8'd168:   begin cos_o = -18'sd72819;  sin_o = 18'sd108982; end
            8'd169:   begin cos_o = -18'sd70123;  sin_o = 18'sd110736; end
            8'd170:   begin cos_o = -18'sd67384;  sin_o = 18'sd112424; end
            8'd171:   begin cos_o = -18'sd64605;  sin_o = 18'sd114044; end
            8'd172:   begin cos_o = -18'sd61786;  sin_o = 18'sd115595; end
            8'd173:   begin cos_o = -18'sd58931;  sin_o = 18'sd117076; end
            8'd174:   begin cos_o = -18'sd56040;  sin_o = 18'sd118487; end
            8'd175:   begin cos_o = -18'sd53115;  sin_o = 18'sd119827; end
            8'd176:   begin cos_o = -18'sd50159;  sin_o = 18'sd121094; end
            8'd177:   begin cos_o = -18'sd47172;  sin_o = 18'sd122289; end
            8'd178:   begin cos_o = -18'sd44156;  sin_o = 18'sd123410; end
            8'd179:   begin cos_o = -18'sd41114;  sin_o = 18'sd124456; end
            8'd180:   begin cos_o = -18'sd38048;  sin_o = 18'sd125428; end
            8'd181:   begin cos_o = -18'sd34958;  sin_o = 18'sd126324; end
            8'd182:   begin cos_o = -18'sd31847;  sin_o = 18'sd127143; end
            8'd183:   begin cos_o = -18'sd28718;  sin_o = 18'sd127887; end
            8'd184:   begin cos_o = -18'sd25570;  sin_o = 18'sd128553; end
            8'd185:   begin cos_o = -18'sd22408;  sin_o = 18'sd129142; end
            8'd186:   begin cos_o = -18'sd19232;  sin_o = 18'sd129653; end
            8'd187:   begin cos_o = -18'sd16044;  sin_o = 18'sd130086; end
            8'd188:   begin cos_o = -18'sd12847;  sin_o = 18'sd130440; end
            8'd189:   begin cos_o = -18'sd9642;  sin_o = 18'sd130716; end
            8'd190:   begin cos_o = -18'sd6431;  sin_o = 18'sd130914; end
            8'd191:   begin cos_o = -18'sd3216;  sin_o = 18'sd131032; end
            8'd192:   begin cos_o = 18'sd0;  sin_o = 18'sd131071; end
            8'd193:   begin cos_o = 18'sd3216;  sin_o = 18'sd131032; end
            8'd194:   begin cos_o = 18'sd6431;  sin_o = 18'sd130914; end
            8'd195:   begin cos_o = 18'sd9642;  sin_o = 18'sd130716; end
            8'd196:   begin cos_o = 18'sd12847;  sin_o = 18'sd130440; end
            8'd197:   begin cos_o = 18'sd16044;  sin_o = 18'sd130086; end
            8'd198:   begin cos_o = 18'sd19232;  sin_o = 18'sd129653; end
            8'd199:   begin cos_o = 18'sd22408;  sin_o = 18'sd129142; end
            8'd200:   begin cos_o = 18'sd25570;  sin_o = 18'sd128553; end
            8'd201:   begin cos_o = 18'sd28718;  sin_o = 18'sd127887; end
            8'd202:   begin cos_o = 18'sd31847;  sin_o = 18'sd127143; end
            8'd203:   begin cos_o = 18'sd34958;  sin_o = 18'sd126324; end
            8'd204:   begin cos_o = 18'sd38048;  sin_o = 18'sd125428; end
            8'd205:   begin cos_o = 18'sd41114;  sin_o = 18'sd124456; end
            8'd206:   begin cos_o = 18'sd44156;  sin_o = 18'sd123410; end
            8'd207:   begin cos_o = 18'sd47172;  sin_o = 18'sd122289; end
            8'd208:   begin cos_o = 18'sd50159;  sin_o = 18'sd121094; end
            8'd209:   begin cos_o = 18'sd53115;  sin_o = 18'sd119827; end
            8'd210:   begin cos_o = 18'sd56040;  sin_o = 18'sd118487; end
            8'd211:   begin cos_o = 18'sd58931;  sin_o = 18'sd117076; end
            8'd212:   begin cos_o = 18'sd61786;  sin_o = 18'sd115595; end
            8'd213:   begin cos_o = 18'sd64605;  sin_o = 18'sd114044; end
            8'd214:   begin cos_o = 18'sd67384;  sin_o = 18'sd112424; end
            8'd215:   begin cos_o = 18'sd70123;  sin_o = 18'sd110736; end
            8'd216:   begin cos_o = 18'sd72819;  sin_o = 18'sd108982; end
            8'd217:   begin cos_o = 18'sd75472;  sin_o = 18'sd107162; end
            8'd218:   begin cos_o = 18'sd78079;  sin_o = 18'sd105278; end
            8'd219:   begin cos_o = 18'sd80639;  sin_o = 18'sd103330; end
            8'd220:   begin cos_o = 18'sd83151;  sin_o = 18'sd101320; end
            8'd221:   begin cos_o = 18'sd85612;  sin_o = 18'sd99248; end
            8'd222:   begin cos_o = 18'sd88022;  sin_o = 18'sd97117; end
            8'd223:   begin cos_o = 18'sd90379;  sin_o = 18'sd94928; end
            8'd224:   begin cos_o = 18'sd92681;  sin_o = 18'sd92681; end
            8'd225:   begin cos_o = 18'sd94928;  sin_o = 18'sd90379; end
            8'd226:   begin cos_o = 18'sd97117;  sin_o = 18'sd88022; end
            8'd227:   begin cos_o = 18'sd99248;  sin_o = 18'sd85612; end
            8'd228:   begin cos_o = 18'sd101320;  sin_o = 18'sd83151; end
            8'd229:   begin cos_o = 18'sd103330;  sin_o = 18'sd80639; end
            8'd230:   begin cos_o = 18'sd105278;  sin_o = 18'sd78079; end
            8'd231:   begin cos_o = 18'sd107162;  sin_o = 18'sd75472; end
            8'd232:   begin cos_o = 18'sd108982;  sin_o = 18'sd72819; end
            8'd233:   begin cos_o = 18'sd110736;  sin_o = 18'sd70123; end
            8'd234:   begin cos_o = 18'sd112424;  sin_o = 18'sd67384; end
            8'd235:   begin cos_o = 18'sd114044;  sin_o = 18'sd64605; end
            8'd236:   begin cos_o = 18'sd115595;  sin_o = 18'sd61786; end
            8'd237:   begin cos_o = 18'sd117076;  sin_o = 18'sd58931; end
            8'd238:   begin cos_o = 18'sd118487;  sin_o = 18'sd56040; end
            8'd239:   begin cos_o = 18'sd119827;  sin_o = 18'sd53115; end
            8'd240:   begin cos_o = 18'sd121094;  sin_o = 18'sd50159; end
            8'd241:   begin cos_o = 18'sd122289;  sin_o = 18'sd47172; end
            8'd242:   begin cos_o = 18'sd123410;  sin_o = 18'sd44156; end
            8'd243:   begin cos_o = 18'sd124456;  sin_o = 18'sd41114; end
            8'd244:   begin cos_o = 18'sd125428;  sin_o = 18'sd38048; end
            8'd245:   begin cos_o = 18'sd126324;  sin_o = 18'sd34958; end
            8'd246:   begin cos_o = 18'sd127143;  sin_o = 18'sd31847; end
            8'd247:   begin cos_o = 18'sd127887;  sin_o = 18'sd28718; end
            8'd248:   begin cos_o = 18'sd128553;  sin_o = 18'sd25570; end
            8'd249:   begin cos_o = 18'sd129142;  sin_o = 18'sd22408; end
            8'd250:   begin cos_o = 18'sd129653;  sin_o = 18'sd19232; end
            8'd251:   begin cos_o = 18'sd130086;  sin_o = 18'sd16044; end
            8'd252:   begin cos_o = 18'sd130440;  sin_o = 18'sd12847; end
            8'd253:   begin cos_o = 18'sd130716;  sin_o = 18'sd9642; end
            8'd254:   begin cos_o = 18'sd130914;  sin_o = 18'sd6431; end
            8'd255:   begin cos_o = 18'sd131032;  sin_o = 18'sd3216; end
        endcase
    end

endmodule
