// removed package "fpga_template_pkg"
module vu_meter_6led (
	clk_i,
	rst_ni,
	sample_stb_i,
	left_sample_i,
	right_sample_i,
	leds_o
);
	reg _sv2v_0;
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:7:13
	parameter [0:0] SELECT_LEFT = 1'b1;
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:8:13
	parameter signed [31:0] DECAY_SHIFT = 11;
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:9:13
	parameter signed [31:0] SCALE_SHIFT = 10;
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:11:13
	parameter [31:0] TH1 = 24'd1000;
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:12:13
	parameter [31:0] TH2 = 24'd3000;
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:13:13
	parameter [31:0] TH3 = 24'd9000;
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:14:13
	parameter [31:0] TH4 = 24'd20000;
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:15:13
	parameter [31:0] TH5 = 24'd40000;
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:16:13
	parameter [31:0] TH6 = 24'd80000;
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:18:13
	parameter signed [31:0] LED_DIV = 540000;
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:20:3
	input wire clk_i;
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:21:3
	input wire rst_ni;
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:22:3
	input wire sample_stb_i;
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:23:3
	input wire signed [23:0] left_sample_i;
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:24:3
	input wire signed [23:0] right_sample_i;
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:25:3
	output reg [5:0] leds_o;
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:28:3
	reg signed [23:0] sample;
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:29:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:29:15
		sample = (SELECT_LEFT ? left_sample_i : right_sample_i);
	end
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:32:3
	reg [23:0] mag;
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:33:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:33:15
		mag = (sample[23] ? ~sample + 1'b1 : sample);
	end
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:36:3
	reg [31:0] level_q;
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:37:3
	always @(posedge clk_i)
		// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:38:5
		if (!rst_ni)
			// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:39:7
			level_q <= 32'd0;
		else if (sample_stb_i)
			// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:42:7
			level_q <= (level_q - (level_q >> DECAY_SHIFT)) + (mag >> SCALE_SHIFT);
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:48:3
	reg [$clog2(LED_DIV) - 1:0] div_q;
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:49:3
	reg tick;
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:50:3
	always @(posedge clk_i)
		// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:51:5
		if (!rst_ni) begin
			// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:52:7
			div_q <= 1'sb0;
			// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:52:20
			tick <= 1'b0;
		end
		else if (div_q == (LED_DIV - 1)) begin
			// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:54:7
			div_q <= 1'sb0;
			// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:54:20
			tick <= 1'b1;
		end
		else begin
			// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:56:7
			div_q <= div_q + 1'b1;
			// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:56:30
			tick <= 1'b0;
		end
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:61:3
	reg [5:0] leds_next;
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:62:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:63:5
		leds_next[0] = level_q > TH1;
		// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:64:5
		leds_next[1] = level_q > TH2;
		// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:65:5
		leds_next[2] = level_q > TH3;
		// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:66:5
		leds_next[3] = level_q > TH4;
		// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:67:5
		leds_next[4] = level_q > TH5;
		// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:68:5
		leds_next[5] = level_q > TH6;
	end
	// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:71:3
	always @(posedge clk_i)
		// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:72:5
		if (!rst_ni)
			// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:72:25
			leds_o <= 6'b000000;
		else if (tick)
			// Trace: /home/tomato-chip/ATKI/digital/sampler/vu_meter_6led.sv:73:25
			leds_o <= leds_next;
	initial _sv2v_0 = 0;
endmodule
